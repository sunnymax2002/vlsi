module soc_top(

);

endmodule